//-------------------------------------------------------------------------------------------------
//  -- ��Ȩ������   : �й���㣨���ţ����޹�˾����ͼ���Ӿ������ֹ�˾, 2010 -2015.
//  -- ���ܼ���     ������.
//  -- ����         : Ӳ������FPGA������
//  -- ģ����       : trigger_active
//  -- �����       : �Ϻ���
//-------------------------------------------------------------------------------------------------
//
//  -- �汾��¼ :
//
//  -- ����         :| �޸�����				:|  �޸�˵��
//-------------------------------------------------------------------------------------------------
//  -- �Ϻ���       :| 2014/12/1 13:25:30	:|  ��ʼ�汾
//-------------------------------------------------------------------------------------------------
//
//  -- ģ������     :��ȡ�����źŵı���
//              1)  : ��С�������źſ����1��ʱ��
//
//              2)  : ����źſ����1��ʱ��
//
//              3)  : ... ...
//
//-------------------------------------------------------------------------------------------------
//���浥λ/����
`timescale 1ns/1ps
//-------------------------------------------------------------------------------------------------

module trigger_active (
	//ϵͳ����
	input			clk					,	//ʱ��72MHz

	//�Ĵ�������
	input			i_trigger_soft		,	//��������
	input	[3:0]	iv_trigger_source	,	//ѡ������Դ��0001-������0010-line0��0100-line2��1000-line3
	input			i_trigger_active	,	//0-�½�����Ч��1��������Ч

	//FPGAģ�齻���ź�
	input			i_din				,	//�����ź�����
	output			o_dout					//�����ź����
	);

	//	ref signals
	reg				triggerl_sel		= 1'b0;	//����Դѡ��
	reg				triggerl_sel_dly	= 1'b0;	//�����źŴ�һ�ģ������ж������źŵı���
	wire			triggerl_sel_rise	;	//�����ر�ʶ
	wire			triggerl_sel_fall	;	//�½��ر�ʶ
	reg				dout_reg			= 1'b0;	//����Ĵ���

	//	ref ARCHITECTURE

	//  -------------------------------------------------------------------------------------
	//	ѡ���ⴥ����������
	//	1.��ѡ������ʱ������Դ�л�Ϊ����
	//	2.��ѡ���ⴥ��ʱ������Դ�л�Ϊ�ⴥ��
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(iv_trigger_source==4'b0001) begin
			triggerl_sel	<= i_trigger_soft;
		end
		else begin
			triggerl_sel	<= i_din;
		end
	end

	//  -------------------------------------------------------------------------------------
	//	�жϱ���
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		triggerl_sel_dly	<= triggerl_sel;
	end
	assign	triggerl_sel_rise	= (triggerl_sel_dly==1'b0 && triggerl_sel==1'b1) ? 1'b1 : 1'b0;
	assign	triggerl_sel_fall	= (triggerl_sel_dly==1'b1 && triggerl_sel==1'b0) ? 1'b1 : 1'b0;

	//  -------------------------------------------------------------------------------------
	//	����ѡ��
	//	0-�½�����Ч��1��������Ч
	//  -------------------------------------------------------------------------------------
	always @ (posedge clk) begin
		if(!i_trigger_active) begin
			dout_reg	<= triggerl_sel_fall;
		end
		else begin
			dout_reg	<= triggerl_sel_rise;
		end
	end
	assign	o_dout	= dout_reg;


endmodule
